-- DIG_OUT.VHD (a peripheral for SCOMP)
-- 2006.10.08
--
-- This device drives 16 digital outputs with data sent from SCOMP.


LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE LPM.LPM_COMPONENTS.ALL;


ENTITY DIG_OUT IS
  PORT(
    RESETN      : IN  STD_LOGIC;
    IO_ADDR     : IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
	 IO_WRITE    : IN  STD_LOGIC;
    IO_DATA     : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
    EXT_WIRES   : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END DIG_OUT;

ARCHITECTURE a OF DIG_OUT IS
  
  SIGNAL CHIP_SELECT : STD_LOGIC;
  
  BEGIN
    CHIP_SELECT <=
      '1' WHEN (IO_ADDR = "00000000001") AND (IO_WRITE = '1')
		ELSE '0';
		
    PROCESS (RESETN, IO_WRITE, CHIP_SELECT)
      BEGIN
        IF (RESETN = '0') THEN
          EXT_WIRES <= x"0000";
        ELSIF (RISING_EDGE(CHIP_SELECT)) THEN
          EXT_WIRES <= IO_DATA;
        END IF;
      END PROCESS;
  END a;

